class transaction;
    integer Data_in;
    logic [3:0] Address;
    logic W_EN;
    logic RST;
    integer Data_out;
endclass