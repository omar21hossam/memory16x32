interface intf;
    logic [31:0]  Data_in;
    logic [3:0] Address;
    logic W_EN;
    logic RST;
    logic CLK;
    logic [31:0]  Data_out;
endinterface