class transaction;
    rand logic [31:0] Data_in;
    randc logic [3:0] Address;
    rand logic W_EN;
    rand logic RST;
    logic [31:0] Data_out;
endclass